
//FUll adder
module fulladder(a,b,c,carry,sum);
input a,b,c;
output sum,carry;
assign sum = a ^ b ^ c;
assign carry = ((a&b)|(b&c)|(c&a));
endmodule

//Half adder
module halfadder(a,b,carry,sum);
input a,b;
output sum,carry;                   
assign sum = a ^ b ;
assign carry = a&b ;
endmodule 

//1-bit flipflop
module flip_flop1(d,q,clk,reset);
input d,clk,reset;
output q;
reg q;
always@(posedge clk)
begin
if(reset==1'b1)
q<=1'b0;
else
q<=d;
end 
endmodule       

//16-bit flip flop
module flip_flop16(d1,q1,clk,reset);
input [15:0] d1;
input clk,reset;
output  [15:0] q1;
reg [15:0] q1;
always@(posedge clk)
begin
if(reset==1'b1)
q1<=16'b0;
else
q1<=d1;
end 
endmodule                  

//multiplier with pipelining            
module mulp(a,b,clk,reset,out);
input [15:0] a,b;
input clk,reset;
output [31:0] out;
wire [15:0]pp0,pp1,pp2,pp3,pp4,pp5,pp6,pp7,pp8,pp9,pp10,pp11,pp12,pp13,pp14,pp15; 
wire [15:0]PP0,PP1,PP2,PP3,PP4,PP5,PP6,PP7,PP8,PP9,PP10,PP11,PP12,PP13,PP14,PP15; 

assign pp0 = {a[15]&b[0],a[14]&b[0],a[13]&b[0],a[12]&b[0],a[11]&b[0],a[10]&b[0],a[9]&b[0],a[8]&b[0],a[7]&b[0],a[6]&b[0],a[5]&b[0],a[4]&b[0],a[3]&b[0],a[2]&b[0],a[1]&b[0],a[0]&b[0]};
assign pp1 = {a[15]&b[1],a[14]&b[1],a[13]&b[1],a[12]&b[1],a[11]&b[1],a[10]&b[1],a[9]&b[1],a[8]&b[1],a[7]&b[1],a[6]&b[1],a[5]&b[1],a[4]&b[1],a[3]&b[1],a[2]&b[1],a[1]&b[1],a[0]&b[1]};
assign pp2 = {a[15]&b[2],a[14]&b[2],a[13]&b[2],a[12]&b[2],a[11]&b[2],a[10]&b[2],a[9]&b[2],a[8]&b[2],a[7]&b[2],a[6]&b[2],a[5]&b[2],a[4]&b[2],a[3]&b[2],a[2]&b[2],a[1]&b[2],a[0]&b[2]};
assign pp3 = {a[15]&b[3],a[14]&b[3],a[13]&b[3],a[12]&b[3],a[11]&b[3],a[10]&b[3],a[9]&b[3],a[8]&b[3],a[7]&b[3],a[6]&b[3],a[5]&b[3],a[4]&b[3],a[3]&b[3],a[2]&b[3],a[1]&b[3],a[0]&b[3]};
assign pp4 = {a[15]&b[4],a[14]&b[4],a[13]&b[4],a[12]&b[4],a[11]&b[4],a[10]&b[4],a[9]&b[4],a[8]&b[4],a[7]&b[4],a[6]&b[4],a[5]&b[4],a[4]&b[4],a[3]&b[4],a[2]&b[4],a[1]&b[4],a[0]&b[4]};
assign pp5 = {a[15]&b[5],a[14]&b[5],a[13]&b[5],a[12]&b[5],a[11]&b[5],a[10]&b[5],a[9]&b[5],a[8]&b[5],a[7]&b[5],a[6]&b[5],a[5]&b[5],a[4]&b[5],a[3]&b[5],a[2]&b[5],a[1]&b[5],a[0]&b[5]};
assign pp6 = {a[15]&b[6],a[14]&b[6],a[13]&b[6],a[12]&b[6],a[11]&b[6],a[10]&b[6],a[9]&b[6],a[8]&b[6],a[7]&b[6],a[6]&b[6],a[5]&b[6],a[4]&b[6],a[3]&b[6],a[2]&b[6],a[1]&b[6],a[0]&b[6]};
assign pp7 = {a[15]&b[7],a[14]&b[7],a[13]&b[7],a[12]&b[7],a[11]&b[7],a[10]&b[7],a[9]&b[7],a[8]&b[7],a[7]&b[7],a[6]&b[7],a[5]&b[7],a[4]&b[7],a[3]&b[7],a[2]&b[7],a[1]&b[7],a[0]&b[7]};
assign pp8 = {a[15]&b[8],a[14]&b[8],a[13]&b[8],a[12]&b[8],a[11]&b[8],a[10]&b[8],a[9]&b[8],a[8]&b[8],a[7]&b[8],a[6]&b[8],a[5]&b[8],a[4]&b[8],a[3]&b[8],a[2]&b[8],a[1]&b[8],a[0]&b[8]};
assign pp9 = {a[15]&b[9],a[14]&b[9],a[13]&b[9],a[12]&b[9],a[11]&b[9],a[10]&b[9],a[9]&b[9],a[8]&b[9],a[7]&b[9],a[6]&b[9],a[5]&b[9],a[4]&b[9],a[3]&b[9],a[2]&b[9],a[1]&b[9],a[0]&b[9]};
assign pp10 = {a[15]&b[10],a[14]&b[10],a[13]&b[10],a[12]&b[10],a[11]&b[10],a[10]&b[10],a[9]&b[10],a[8]&b[10],a[7]&b[10],a[6]&b[10],a[5]&b[10],a[4]&b[10],a[3]&b[10],a[2]&b[10],a[1]&b[10],a[0]&b[10]};
assign pp11 = {a[15]&b[11],a[14]&b[11],a[13]&b[11],a[12]&b[11],a[11]&b[11],a[10]&b[11],a[9]&b[11],a[8]&b[11],a[7]&b[11],a[6]&b[11],a[5]&b[11],a[4]&b[11],a[3]&b[11],a[2]&b[11],a[1]&b[11],a[0]&b[11]};
assign pp12 = {a[15]&b[12],a[14]&b[12],a[13]&b[12],a[12]&b[12],a[11]&b[12],a[10]&b[12],a[9]&b[12],a[8]&b[12],a[7]&b[12],a[6]&b[12],a[5]&b[12],a[4]&b[12],a[3]&b[12],a[2]&b[12],a[1]&b[12],a[0]&b[12]};
assign pp13 = {a[15]&b[13],a[14]&b[13],a[13]&b[13],a[12]&b[13],a[11]&b[13],a[10]&b[13],a[9]&b[13],a[8]&b[13],a[7]&b[13],a[6]&b[13],a[5]&b[13],a[4]&b[13],a[3]&b[13],a[2]&b[13],a[1]&b[13],a[0]&b[13]};
assign pp14 = {a[15]&b[14],a[14]&b[14],a[13]&b[14],a[12]&b[14],a[11]&b[14],a[10]&b[14],a[9]&b[14],a[8]&b[14],a[7]&b[14],a[6]&b[14],a[5]&b[14],a[4]&b[14],a[3]&b[14],a[2]&b[14],a[1]&b[14],a[0]&b[14]};
assign pp15 = {a[15]&b[15],a[14]&b[15],a[13]&b[15],a[12]&b[15],a[11]&b[15],a[10]&b[15],a[9]&b[15],a[8]&b[15],a[7]&b[15],a[6]&b[15],a[5]&b[15],a[4]&b[15],a[3]&b[15],a[2]&b[15],a[1]&b[15],a[0]&b[15]};      
   
wire [15:0]a1PP2,a1PP3,a1PP4,a1PP5,a1PP6,a1PP7,a1PP8,a1PP9,a1PP10,a1PP11,a1PP12,a1PP13,a1PP14,a1PP15;
wire [15:0]b2PP3,b2PP4,b2PP5,b2PP6,b2PP7,b2PP8,b2PP9,b2PP10,b2PP11,b2PP12,b2PP13,b2PP14,b2PP15;    
wire [15:0]c3PP4,c3PP5,c3PP6,c3PP7,c3PP8,c3PP9,c3PP10,c3PP11,c3PP12,c3PP13,c3PP14,c3PP15;         
wire [15:0]d4PP5,d4PP6,d4PP7,d4PP8,d4PP9,d4PP10,d4PP11,d4PP12,d4PP13,d4PP14,d4PP15;              
wire [15:0]e5PP6,e5PP7,e5PP8,e5PP9,e5PP10,e5PP11,e5PP12,e5PP13,e5PP14,e5PP15;                   
wire [15:0]f6PP7,f6PP8,f6PP9,f6PP10,f6PP11,f6PP12,f6PP13,f6PP14,f6PP15;                        
wire [15:0]g7PP8,g7PP9,g7PP10,g7PP11,g7PP12,g7PP13,g7PP14,g7PP15;                             
wire [15:0]h8PP9,h8PP10,h8PP11,h8PP12,h8PP13,h8PP14,h8PP15;                                  
wire [15:0]i9PP10,i9PP11,i9PP12,i9PP13,i9PP14,i9PP15;                                       
wire [15:0]j10PP11,j10PP12,j10PP13,j10PP14,j10PP15;                                        
wire [15:0]k11PP12,k11PP13,k11PP14,k11PP15;                                               
wire [15:0]l12PP13,l12PP14,l12PP15;                                                      
wire [15:0]m13PP14,m13PP15;                                                             
wire [15:0]n14PP15; 

flip_flop16 mod1400(pp0,PP0,clk,reset);
flip_flop16 mod1300(pp1,PP1,clk,reset);
flip_flop16 mod1301(pp2,PP2,clk,reset);
flip_flop16 mod1302(pp3,PP3,clk,reset);
flip_flop16 mod1303(pp4,PP4,clk,reset);
flip_flop16 mod1304(pp5,PP5,clk,reset);
flip_flop16 mod1305(pp6,PP6,clk,reset);
flip_flop16 mod1306(pp7,PP7,clk,reset);
flip_flop16 mod1307(pp8,PP8,clk,reset);
flip_flop16 mod1308(pp9,PP9,clk,reset);
flip_flop16 mod1309(pp10,PP10,clk,reset);
flip_flop16 mod1310(pp11,PP11,clk,reset);
flip_flop16 mod1311(pp12,PP12,clk,reset);
flip_flop16 mod1312(pp13,PP13,clk,reset);
flip_flop16 mod1313(pp14,PP14,clk,reset);
flip_flop16 mod1314(pp15,PP15,clk,reset);
//FOR STAGE - 1
assign p0 = PP0[0];
halfadder mod0(PP0[1],PP1[0],carry1,p1);
fulladder mod1(PP0[2],PP1[1],PP2[0],carry2,sum1);
fulladder mod2(PP0[3],PP1[2],PP2[1],carry3,sum2);
fulladder mod3(PP0[4],PP1[3],PP2[2],carry4,sum3);
fulladder mod4(PP0[5],PP1[4],PP2[3],carry5,sum4);
fulladder mod5(PP0[6],PP1[5],PP2[4],carry6,sum5);
fulladder mod6(PP0[7],PP1[6],PP2[5],carry7,sum6);
fulladder mod7(PP0[8],PP1[7],PP2[6],carry8,sum7);
fulladder mod8(PP0[9],PP1[8],PP2[7],carry9,sum8);
fulladder mod9(PP0[10],PP1[9],PP2[8],carry10,sum9);
fulladder mod10(PP0[11],PP1[10],PP2[9],carry11,sum10);
fulladder mod11(PP0[12],PP1[11],PP2[10],carry12,sum11);
fulladder mod12(PP0[13],PP1[12],PP2[11],carry13,sum12);
fulladder mod13(PP0[14],PP1[13],PP2[12],carry14,sum13);
fulladder mod14(PP0[15],PP1[14],PP2[13],carry15,sum14);                                                                       
//FOR STAGE - 1 PIPELINE 
flip_flop1 mod241(p0,p01,clk,reset); 
flip_flop1 mod242(p1,p11,clk,reset); 
flip_flop1 mod243(carry1,qcarry1,clk,reset); 
flip_flop1 mod244(carry2,qcarry2,clk,reset);
flip_flop1 mod245(carry3,qcarry3,clk,reset);
flip_flop1 mod246(carry4,qcarry4,clk,reset);
flip_flop1 mod247(carry5,qcarry5,clk,reset);
flip_flop1 mod248(carry6,qcarry6,clk,reset);
flip_flop1 mod249(carry7,qcarry7,clk,reset); 
flip_flop1 mod250(carry8,qcarry8,clk,reset); 
flip_flop1 mod251(carry9,qcarry9,clk,reset); 
flip_flop1 mod252(carry10,qcarry10,clk,reset);
flip_flop1 mod253(carry11,qcarry11,clk,reset);
flip_flop1 mod254(carry12,qcarry12,clk,reset);
flip_flop1 mod255(carry13,qcarry13,clk,reset);     
flip_flop1 mod256(carry14,qcarry14,clk,reset);
flip_flop1 mod257(carry15,qcarry15,clk,reset); 

flip_flop1  mod258(sum1,qsum1,clk,reset); 
flip_flop1  mod259(sum2,qsum2,clk,reset);
flip_flop1  mod260(sum3,qsum3,clk,reset);
flip_flop1  mod261(sum4,qsum4,clk,reset);
flip_flop1  mod262(sum5,qsum5,clk,reset);
flip_flop1  mod263(sum6,qsum6,clk,reset); 
flip_flop1  mod264(sum7,qsum7,clk,reset); 
flip_flop1  mod265(sum8,qsum8,clk,reset);
flip_flop1  mod266(sum9,qsum9,clk,reset);
flip_flop1  mod267(sum10,qsum10,clk,reset);
flip_flop1  mod268(sum11,qsum11,clk,reset);
flip_flop1  mod269(sum12,qsum12,clk,reset);
flip_flop1  mod270(sum13,qsum13,clk,reset);
flip_flop1  mod271(sum14,qsum14,clk,reset); 

flip_flop1 mod1000(PP1[15],a1PP1,clk,reset);
flip_flop16 mod1001(PP2,a1PP2,clk,reset);
flip_flop16 mod1002(PP3,a1PP3,clk,reset);
flip_flop16 mod1003(PP4,a1PP4,clk,reset);
flip_flop16 mod1004(PP5,a1PP5,clk,reset);
flip_flop16 mod1005(PP6,a1PP6,clk,reset);
flip_flop16 mod1006(PP7,a1PP7,clk,reset);
flip_flop16 mod1007(PP8,a1PP8,clk,reset);
flip_flop16 mod1008(PP9,a1PP9,clk,reset);
flip_flop16 mod1009(PP10,a1PP10,clk,reset);
flip_flop16 mod1010(PP11,a1PP11,clk,reset);
flip_flop16 mod1011(PP12,a1PP12,clk,reset);
flip_flop16 mod1012(PP13,a1PP13,clk,reset);
flip_flop16 mod1013(PP14,a1PP14,clk,reset);
flip_flop16 mod1014(PP15,a1PP15,clk,reset);
//FOR STAGE - 2   
halfadder mod15(qsum1,qcarry1,carry16,p2);
fulladder mod16(qsum2,qcarry2,a1PP3[0],carry17,sum15);  
fulladder mod17(qsum3,qcarry3,a1PP3[1],carry18,sum16);                                            
fulladder mod18(qsum4,qcarry4,a1PP3[2],carry19,sum17);
fulladder mod19(qsum5,qcarry5,a1PP3[3],carry20,sum18);
fulladder mod20(qsum6,qcarry6,a1PP3[4],carry21,sum19);
fulladder mod21(qsum7,qcarry7,a1PP3[5],carry22,sum20);
fulladder mod22(qsum8,qcarry8,a1PP3[6],carry23,sum21);
fulladder mod23(qsum9,qcarry9,a1PP3[7],carry24,sum22);
fulladder mod24(qsum10,qcarry10,a1PP3[8],carry25,sum23);
fulladder mod25(qsum11,qcarry11,a1PP3[9],carry26,sum24);
fulladder mod26(qsum12,qcarry12,a1PP3[10],carry27,sum25);
fulladder mod27(qsum13,qcarry13,a1PP3[11],carry28,sum26);
fulladder mod28(qsum14,qcarry14,a1PP3[12],carry29,sum27);
fulladder mod29(a1PP1,a1PP2[14],qcarry15,carry30,sum28);
//FOR STAGE - 2 PIPELINE 
flip_flop1  mod272(p01,p02,clk,reset); 
flip_flop1  mod273(p11,p12,clk,reset);
flip_flop1  mod274(p2,p21,clk,reset); 
flip_flop1  mod275(carry16,qcarry16,clk,reset); 
flip_flop1  mod276(carry17,qcarry17,clk,reset);
flip_flop1  mod277(carry18,qcarry18,clk,reset);
flip_flop1  mod278(carry19,qcarry19,clk,reset);
flip_flop1  mod279(carry20,qcarry20,clk,reset);
flip_flop1  mod280(carry21,qcarry21,clk,reset);
flip_flop1  mod281(carry22,qcarry22,clk,reset); 
flip_flop1  mod282(carry23,qcarry23,clk,reset); 
flip_flop1  mod283(carry24,qcarry24,clk,reset); 
flip_flop1  mod284(carry25,qcarry25,clk,reset);
flip_flop1  mod285(carry26,qcarry26,clk,reset);
flip_flop1  mod286(carry27,qcarry27,clk,reset);
flip_flop1  mod287(carry28,qcarry28,clk,reset);     
flip_flop1  mod288(carry29,qcarry29,clk,reset);
flip_flop1  mod289(carry30,qcarry30,clk,reset); 
          
flip_flop1  mod290(sum15,qsum15,clk,reset);
flip_flop1  mod291(sum16,qsum16,clk,reset);
flip_flop1  mod292(sum17,qsum17,clk,reset);
flip_flop1  mod293(sum18,qsum18,clk,reset);
flip_flop1  mod294(sum19,qsum19,clk,reset);
flip_flop1  mod295(sum20,qsum20,clk,reset);
flip_flop1  mod296(sum21,qsum21,clk,reset);
flip_flop1  mod297(sum22,qsum22,clk,reset);
flip_flop1  mod298(sum23,qsum23,clk,reset);
flip_flop1  mod299(sum24,qsum24,clk,reset);
flip_flop1  mod300(sum25,qsum25,clk,reset);
flip_flop1  mod301(sum26,qsum26,clk,reset);
flip_flop1  mod302(sum27,qsum27,clk,reset);
flip_flop1  mod303(sum28,qsum28,clk,reset); 

flip_flop1 mod1015(a1PP2[15],b2PP2,clk,reset);
flip_flop16 mod1016(a1PP3,b2PP3,clk,reset);
flip_flop16 mod1017(a1PP4,b2PP4,clk,reset);
flip_flop16 mod1018(a1PP5,b2PP5,clk,reset);
flip_flop16 mod1019(a1PP6,b2PP6,clk,reset);
flip_flop16 mod1020(a1PP7,b2PP7,clk,reset);
flip_flop16 mod1021(a1PP8,b2PP8,clk,reset);
flip_flop16 mod1022(a1PP9,b2PP9,clk,reset);
flip_flop16 mod1023(a1PP10,b2PP10,clk,reset);
flip_flop16 mod1024(a1PP11,b2PP11,clk,reset);
flip_flop16 mod1025(a1PP12,b2PP12,clk,reset);
flip_flop16 mod1026(a1PP13,b2PP13,clk,reset);
flip_flop16 mod1027(a1PP14,b2PP14,clk,reset);
flip_flop16 mod1028(a1PP15,b2PP15,clk,reset);
//FOR STAGE - 3
halfadder mod30(qsum15,qcarry16,carry31,p3);
fulladder mod31(qsum16,qcarry17,b2PP4[0],carry32,sum29);  
fulladder mod32(qsum17,qcarry18,b2PP4[1],carry33,sum30);
fulladder mod33(qsum18,qcarry19,b2PP4[2],carry34,sum31);
fulladder mod34(qsum19,qcarry20,b2PP4[3],carry35,sum32);
fulladder mod35(qsum20,qcarry21,b2PP4[4],carry36,sum33);
fulladder mod36(qsum21,qcarry22,b2PP4[5],carry37,sum34);
fulladder mod37(qsum22,qcarry23,b2PP4[6],carry38,sum35);
fulladder mod38(qsum23,qcarry24,b2PP4[7],carry39,sum36);
fulladder mod39(qsum24,qcarry25,b2PP4[8],carry40,sum37);
fulladder mod40(qsum25,qcarry26,b2PP4[9],carry41,sum38);
fulladder mod41(qsum26,qcarry27,b2PP4[10],carry42,sum39);
fulladder mod42(qsum27,qcarry28,b2PP4[11],carry43,sum40);
fulladder mod43(qsum28,qcarry29,b2PP3[13],carry44,sum41);
fulladder mod44(b2PP2,b2PP3[14],qcarry30,carry45,sum42);
//FOR STAGE - 3 PIPELINE 
flip_flop1  mod304(p02,p03,clk,reset); 
flip_flop1  mod305(p12,p13,clk,reset);
flip_flop1  mod306(p21,p22,clk,reset);
flip_flop1  mod307(p3,p31,clk,reset);
flip_flop1  mod308(carry31,qcarry31,clk,reset); 
flip_flop1  mod309(carry32,qcarry32,clk,reset);
flip_flop1  mod310(carry33,qcarry33,clk,reset);
flip_flop1  mod311(carry34,qcarry34,clk,reset);
flip_flop1  mod312(carry35,qcarry35,clk,reset);
flip_flop1  mod313(carry36,qcarry36,clk,reset);
flip_flop1  mod314(carry37,qcarry37,clk,reset); 
flip_flop1  mod315(carry38,qcarry38,clk,reset); 
flip_flop1  mod316(carry39,qcarry39,clk,reset); 
flip_flop1  mod317(carry40,qcarry40,clk,reset);
flip_flop1  mod318(carry41,qcarry41,clk,reset);
flip_flop1  mod319(carry42,qcarry42,clk,reset);
flip_flop1  mod320(carry43,qcarry43,clk,reset);     
flip_flop1  mod321(carry44,qcarry44,clk,reset);
flip_flop1  mod322(carry45,qcarry45,clk,reset); 
         
flip_flop1  mod323(sum29,qsum29,clk,reset);
flip_flop1  mod324(sum30,qsum30,clk,reset);
flip_flop1  mod325(sum31,qsum31,clk,reset);
flip_flop1  mod326(sum32,qsum32,clk,reset);
flip_flop1  mod327(sum33,qsum33,clk,reset);
flip_flop1  mod328(sum34,qsum34,clk,reset);
flip_flop1  mod329(sum35,qsum35,clk,reset);
flip_flop1  mod330(sum36,qsum36,clk,reset);
flip_flop1  mod331(sum37,qsum37,clk,reset);
flip_flop1  mod332(sum38,qsum38,clk,reset);
flip_flop1  mod333(sum39,qsum39,clk,reset);
flip_flop1  mod334(sum40,qsum40,clk,reset);
flip_flop1  mod335(sum41,qsum41,clk,reset);
flip_flop1  mod336(sum42,qsum42,clk,reset);

flip_flop1 mod1029(b2PP3[15],c3PP3,clk,reset);
flip_flop16 mod1031(b2PP4,c3PP4,clk,reset);
flip_flop16 mod1032(b2PP5,c3PP5,clk,reset);
flip_flop16 mod1033(b2PP6,c3PP6,clk,reset);
flip_flop16 mod1034(b2PP7,c3PP7,clk,reset);
flip_flop16 mod1035(b2PP8,c3PP8,clk,reset);
flip_flop16 mod1036(b2PP9,c3PP9,clk,reset);
flip_flop16 mod1037(b2PP10,c3PP10,clk,reset);
flip_flop16 mod1038(b2PP11,c3PP11,clk,reset);
flip_flop16 mod1039(b2PP12,c3PP12,clk,reset);
flip_flop16 mod1040(b2PP13,c3PP13,clk,reset);
flip_flop16 mod1041(b2PP14,c3PP14,clk,reset);
flip_flop16 mod1042(b2PP15,c3PP15,clk,reset);
//FOR STAGE - 4
halfadder mod45(qsum29,qcarry31,carry46,p4);
fulladder mod46(qsum30,qcarry32,c3PP5[0],carry47,sum43);  
fulladder mod47(qsum31,qcarry33,c3PP5[1],carry48,sum44);
fulladder mod48(qsum32,qcarry34,c3PP5[2],carry49,sum45);
fulladder mod49(qsum33,qcarry35,c3PP5[3],carry50,sum46);
fulladder mod50(qsum34,qcarry36,c3PP5[4],carry51,sum47);
fulladder mod51(qsum35,qcarry37,c3PP5[5],carry52,sum48);
fulladder mod52(qsum36,qcarry38,c3PP5[6],carry53,sum49);
fulladder mod53(qsum37,qcarry39,c3PP5[7],carry54,sum50);
fulladder mod54(qsum38,qcarry40,c3PP5[8],carry55,sum51);
fulladder mod55(qsum39,qcarry41,c3PP5[9],carry56,sum52);
fulladder mod56(qsum40,qcarry42,c3PP5[10],carry57,sum53);
fulladder mod57(qsum41,qcarry43,c3PP4[12],carry58,sum54);
fulladder mod58(qsum42,qcarry44,c3PP4[13],carry59,sum55);
fulladder mod59(c3PP3,c3PP4[14],qcarry45,carry60,sum56);
//FOR STAGE - 4 PIPELINE 
flip_flop1  mod337(p03,p04,clk,reset); 
flip_flop1  mod338(p13,p14,clk,reset);
flip_flop1  mod339(p22,p23,clk,reset);
flip_flop1  mod340(p31,p32,clk,reset);
flip_flop1  mod341(p4,p41,clk,reset);
flip_flop1  mod342(carry46,qcarry46,clk,reset); 
flip_flop1  mod343(carry47,qcarry47,clk,reset);
flip_flop1  mod344(carry48,qcarry48,clk,reset);
flip_flop1  mod345(carry49,qcarry49,clk,reset);
flip_flop1  mod346(carry50,qcarry50,clk,reset);
flip_flop1  mod347(carry51,qcarry51,clk,reset);
flip_flop1  mod348(carry52,qcarry52,clk,reset); 
flip_flop1  mod349(carry53,qcarry53,clk,reset); 
flip_flop1  mod350(carry54,qcarry54,clk,reset); 
flip_flop1  mod351(carry55,qcarry55,clk,reset);
flip_flop1  mod352(carry56,qcarry56,clk,reset);
flip_flop1  mod353(carry57,qcarry57,clk,reset);
flip_flop1  mod354(carry58,qcarry58,clk,reset);     
flip_flop1  mod355(carry59,qcarry59,clk,reset);
flip_flop1  mod356(carry60,qcarry60,clk,reset); 
         
flip_flop1  mod357(sum43,qsum43,clk,reset);
flip_flop1  mod358(sum44,qsum44,clk,reset);
flip_flop1  mod359(sum45,qsum45,clk,reset);
flip_flop1  mod360(sum46,qsum46,clk,reset);
flip_flop1  mod361(sum47,qsum47,clk,reset);
flip_flop1  mod362(sum48,qsum48,clk,reset);
flip_flop1  mod363(sum49,qsum49,clk,reset);
flip_flop1  mod364(sum50,qsum50,clk,reset);
flip_flop1  mod365(sum51,qsum51,clk,reset);
flip_flop1  mod366(sum52,qsum52,clk,reset);
flip_flop1  mod367(sum53,qsum53,clk,reset);
flip_flop1  mod368(sum54,qsum54,clk,reset);
flip_flop1  mod369(sum55,qsum55,clk,reset);
flip_flop1  mod370(sum56,qsum56,clk,reset);  
  
flip_flop1 mod1043(c3PP4[15],d4PP4,clk,reset);
flip_flop16  mod1044(c3PP5,d4PP5,clk,reset);
flip_flop16  mod1045(c3PP6,d4PP6,clk,reset);
flip_flop16  mod1046(c3PP7,d4PP7,clk,reset);
flip_flop16  mod1047(c3PP8,d4PP8,clk,reset);
flip_flop16  mod1048(c3PP9,d4PP9,clk,reset);
flip_flop16  mod1049(c3PP10,d4PP10,clk,reset);
flip_flop16  mod1050(c3PP11,d4PP11,clk,reset);
flip_flop16  mod1051(c3PP12,d4PP12,clk,reset);
flip_flop16  mod1052(c3PP13,d4PP13,clk,reset);
flip_flop16  mod1053(c3PP14,d4PP14,clk,reset);
flip_flop16  mod1054(c3PP15,d4PP15,clk,reset);
//FOR STAGE - 5
halfadder mod60(qsum43,qcarry46,carry61,p5);
fulladder mod61(qsum44,qcarry47,d4PP6[0],carry62,sum57);  
fulladder mod62(qsum45,qcarry48,d4PP6[1],carry63,sum58);
fulladder mod63(qsum46,qcarry49,d4PP6[2],carry64,sum59);
fulladder mod64(qsum47,qcarry50,d4PP6[3],carry65,sum60);
fulladder mod65(qsum48,qcarry51,d4PP6[4],carry66,sum61);
fulladder mod66(qsum49,qcarry52,d4PP6[5],carry67,sum62);
fulladder mod67(qsum50,qcarry53,d4PP6[6],carry68,sum63);
fulladder mod68(qsum51,qcarry54,d4PP6[7],carry69,sum64);
fulladder mod69(qsum52,qcarry55,d4PP6[8],carry70,sum65);
fulladder mod70(qsum53,qcarry56,d4PP6[9],carry71,sum66);
fulladder mod71(qsum54,qcarry57,d4PP5[11],carry72,sum67);
fulladder mod72(qsum55,qcarry58,d4PP5[12],carry73,sum68);
fulladder mod73(qsum56,qcarry59,d4PP5[13],carry74,sum69);
fulladder mod74(d4PP4,d4PP5[14],qcarry60,carry75,sum70);
//FOR STAGE - 5 PIPELINE 
flip_flop1  mod371(p04,p05,clk,reset); 
flip_flop1  mod372(p14,p15,clk,reset);
flip_flop1  mod373(p23,p24,clk,reset);
flip_flop1  mod374(p32,p33,clk,reset);
flip_flop1  mod375(p41,p42,clk,reset);
flip_flop1  mod376(p5,p51,clk,reset);
flip_flop1  mod377(carry61,qcarry61,clk,reset); 
flip_flop1  mod378(carry62,qcarry62,clk,reset);
flip_flop1  mod379(carry63,qcarry63,clk,reset);
flip_flop1  mod380(carry64,qcarry64,clk,reset);
flip_flop1  mod381(carry65,qcarry65,clk,reset);
flip_flop1  mod382(carry66,qcarry66,clk,reset);
flip_flop1  mod383(carry67,qcarry67,clk,reset); 
flip_flop1  mod384(carry68,qcarry68,clk,reset); 
flip_flop1  mod385(carry69,qcarry69,clk,reset); 
flip_flop1  mod386(carry70,qcarry70,clk,reset);
flip_flop1  mod387(carry71,qcarry71,clk,reset);
flip_flop1  mod388(carry72,qcarry72,clk,reset);
flip_flop1  mod389(carry73,qcarry73,clk,reset);     
flip_flop1  mod390(carry74,qcarry74,clk,reset);
flip_flop1  mod391(carry75,qcarry75,clk,reset); 
         
flip_flop1  mod392(sum57,qsum57,clk,reset);
flip_flop1  mod393(sum58,qsum58,clk,reset);
flip_flop1  mod394(sum59,qsum59,clk,reset);
flip_flop1  mod395(sum60,qsum60,clk,reset);
flip_flop1  mod396(sum61,qsum61,clk,reset);
flip_flop1  mod397(sum62,qsum62,clk,reset);
flip_flop1  mod398(sum63,qsum63,clk,reset);
flip_flop1  mod399(sum64,qsum64,clk,reset);
flip_flop1  mod400(sum65,qsum65,clk,reset);
flip_flop1  mod401(sum66,qsum66,clk,reset);
flip_flop1  mod402(sum67,qsum67,clk,reset);
flip_flop1  mod403(sum68,qsum68,clk,reset);
flip_flop1  mod404(sum69,qsum69,clk,reset);
flip_flop1  mod405(sum70,qsum70,clk,reset);          
         
flip_flop1 mod1055(d4PP5[15],e5PP5,clk,reset);
flip_flop16  mod1056(d4PP6,e5PP6,clk,reset);
flip_flop16  mod1057(d4PP7,e5PP7,clk,reset);
flip_flop16  mod1058(d4PP8,e5PP8,clk,reset);
flip_flop16  mod1059(d4PP9,e5PP9,clk,reset);
flip_flop16  mod1060(d4PP10,e5PP10,clk,reset);
flip_flop16  mod1061(d4PP11,e5PP11,clk,reset);
flip_flop16  mod1062(d4PP12,e5PP12,clk,reset);
flip_flop16  mod1063(d4PP13,e5PP13,clk,reset);
flip_flop16  mod1064(d4PP14,e5PP14,clk,reset);
flip_flop16  mod1065(d4PP15,e5PP15,clk,reset);
//FOR STAGE - 6 
halfadder mod75(qsum57,qcarry61,carry76,p6);
fulladder mod76(qsum58,qcarry62,e5PP7[0],carry77,sum71);  
fulladder mod77(qsum59,qcarry63,e5PP7[1],carry78,sum72);
fulladder mod78(qsum60,qcarry64,e5PP7[2],carry79,sum73);
fulladder mod79(qsum61,qcarry65,e5PP7[3],carry80,sum74);
fulladder mod80(qsum62,qcarry66,e5PP7[4],carry81,sum75);
fulladder mod81(qsum63,qcarry67,e5PP7[5],carry82,sum76);
fulladder mod82(qsum64,qcarry68,e5PP7[6],carry83,sum77);
fulladder mod83(qsum65,qcarry69,e5PP7[7],carry84,sum78);
fulladder mod84(qsum66,qcarry70,e5PP7[8],carry85,sum79);
fulladder mod85(qsum67,qcarry71,e5PP6[10],carry86,sum80);
fulladder mod86(qsum68,qcarry72,e5PP6[11],carry87,sum81);
fulladder mod87(qsum69,qcarry73,e5PP6[12],carry88,sum82);
fulladder mod88(qsum70,qcarry74,e5PP6[13],carry89,sum83);
fulladder mod89(e5PP5,e5PP6[14],qcarry75,carry90,sum84);
//FOR STAGE - 6 PIPELINE 
flip_flop1  mod406(p05,p06,clk,reset); 
flip_flop1  mod407(p15,p16,clk,reset);
flip_flop1  mod408(p24,p25,clk,reset);
flip_flop1  mod409(p33,p34,clk,reset);
flip_flop1  mod410(p42,p43,clk,reset);
flip_flop1  mod411(p51,p52,clk,reset);
flip_flop1  mod412(p6,p61,clk,reset);
flip_flop1  mod413(carry76,qcarry76,clk,reset); 
flip_flop1  mod414(carry77,qcarry77,clk,reset);
flip_flop1  mod415(carry78,qcarry78,clk,reset);
flip_flop1  mod416(carry79,qcarry79,clk,reset);
flip_flop1  mod417(carry80,qcarry80,clk,reset);
flip_flop1  mod418(carry81,qcarry81,clk,reset);
flip_flop1  mod419(carry82,qcarry82,clk,reset); 
flip_flop1  mod420(carry83,qcarry83,clk,reset); 
flip_flop1  mod421(carry84,qcarry84,clk,reset); 
flip_flop1  mod422(carry85,qcarry85,clk,reset);
flip_flop1  mod423(carry86,qcarry86,clk,reset);
flip_flop1  mod424(carry87,qcarry87,clk,reset);
flip_flop1  mod425(carry88,qcarry88,clk,reset);     
flip_flop1  mod426(carry89,qcarry89,clk,reset);
flip_flop1  mod427(carry90,qcarry90,clk,reset); 
         
flip_flop1  mod428(sum71,qsum71,clk,reset);
flip_flop1  mod429(sum72,qsum72,clk,reset);
flip_flop1  mod430(sum73,qsum73,clk,reset);
flip_flop1  mod431(sum74,qsum74,clk,reset);
flip_flop1  mod432(sum75,qsum75,clk,reset);
flip_flop1  mod433(sum76,qsum76,clk,reset);
flip_flop1  mod434(sum77,qsum77,clk,reset);
flip_flop1  mod435(sum78,qsum78,clk,reset);
flip_flop1  mod436(sum79,qsum79,clk,reset);
flip_flop1  mod437(sum80,qsum80,clk,reset);
flip_flop1  mod438(sum81,qsum81,clk,reset);
flip_flop1  mod439(sum82,qsum82,clk,reset);
flip_flop1  mod440(sum83,qsum83,clk,reset);
flip_flop1  mod441(sum84,qsum84,clk,reset);

flip_flop1 mod1066(e5PP6[15],f6PP6,clk,reset);
flip_flop16  mod1067(e5PP7,f6PP7,clk,reset);
flip_flop16  mod1068(e5PP8,f6PP8,clk,reset);
flip_flop16  mod1069(e5PP9,f6PP9,clk,reset);
flip_flop16  mod1070(e5PP10,f6PP10,clk,reset);
flip_flop16  mod1071(e5PP11,f6PP11,clk,reset);
flip_flop16  mod1072(e5PP12,f6PP12,clk,reset);
flip_flop16  mod1073(e5PP13,f6PP13,clk,reset);
flip_flop16  mod1074(e5PP14,f6PP14,clk,reset);
flip_flop16  mod1075(e5PP15,f6PP15,clk,reset);
//FOR STAGE - 7
halfadder mod90(qsum71,qcarry76,carry91,p7);
fulladder mod91(qsum72,qcarry77,f6PP8[0],carry92,sum85);  
fulladder mod92(qsum73,qcarry78,f6PP8[1],carry93,sum86);
fulladder mod93(qsum74,qcarry79,f6PP8[2],carry94,sum87);
fulladder mod94(qsum75,qcarry80,f6PP8[3],carry95,sum88);
fulladder mod95(qsum76,qcarry81,f6PP8[4],carry96,sum89);
fulladder mod96(qsum77,qcarry82,f6PP8[5],carry97,sum90);
fulladder mod97(qsum78,qcarry83,f6PP8[6],carry98,sum91);
fulladder mod98(qsum79,qcarry84,f6PP8[7],carry99,sum92);
fulladder mod99(qsum80,qcarry85,f6PP7[9],carry100,sum93);
fulladder mod100(qsum81,qcarry86,f6PP7[10],carry101,sum94);
fulladder mod101(qsum82,qcarry87,f6PP7[11],carry102,sum95);
fulladder mod102(qsum83,qcarry88,f6PP7[12],carry103,sum96);
fulladder mod103(qsum84,qcarry89,f6PP7[13],carry104,sum97);
fulladder mod104(f6PP6,f6PP7[14],qcarry90,carry105,sum98);
//FOR STAGE - 7 PIPELINE 
flip_flop1  mod442(p06,p07,clk,reset); 
flip_flop1  mod443(p16,p17,clk,reset);
flip_flop1  mod444(p25,p26,clk,reset);
flip_flop1  mod445(p34,p35,clk,reset);
flip_flop1  mod446(p43,p44,clk,reset);
flip_flop1  mod447(p52,p53,clk,reset);
flip_flop1  mod448(p61,p62,clk,reset);
flip_flop1  mod449(p7,p71,clk,reset);
flip_flop1  mod450(carry91,qcarry91,clk,reset); 
flip_flop1  mod451(carry92,qcarry92,clk,reset);
flip_flop1  mod452(carry93,qcarry93,clk,reset);
flip_flop1  mod453(carry94,qcarry94,clk,reset);
flip_flop1  mod454(carry95,qcarry95,clk,reset);
flip_flop1  mod455(carry96,qcarry96,clk,reset);
flip_flop1  mod456(carry97,qcarry97,clk,reset); 
flip_flop1  mod457(carry98,qcarry98,clk,reset); 
flip_flop1  mod458(carry99,qcarry99,clk,reset); 
flip_flop1  mod459(carry100,qcarry100,clk,reset);
flip_flop1  mod460(carry101,qcarry101,clk,reset);
flip_flop1  mod461(carry102,qcarry102,clk,reset);
flip_flop1  mod462(carry103,qcarry103,clk,reset);     
flip_flop1  mod463(carry104,qcarry104,clk,reset);
flip_flop1  mod464(carry105,qcarry105,clk,reset); 
         
flip_flop1  mod465(sum85,qsum85,clk,reset);
flip_flop1  mod466(sum86,qsum86,clk,reset);
flip_flop1  mod467(sum87,qsum87,clk,reset);
flip_flop1  mod468(sum88,qsum88,clk,reset);
flip_flop1  mod469(sum89,qsum89,clk,reset);
flip_flop1  mod470(sum90,qsum90,clk,reset);
flip_flop1  mod471(sum91,qsum91,clk,reset);
flip_flop1  mod472(sum92,qsum92,clk,reset);
flip_flop1  mod473(sum93,qsum93,clk,reset);
flip_flop1  mod474(sum94,qsum94,clk,reset);
flip_flop1  mod475(sum95,qsum95,clk,reset);
flip_flop1  mod476(sum96,qsum96,clk,reset);
flip_flop1  mod477(sum97,qsum97,clk,reset);
flip_flop1  mod478(sum98,qsum98,clk,reset);

flip_flop1 mod1076(f6PP7[15],g7PP7,clk,reset);
flip_flop16  mod1077(f6PP8,g7PP8,clk,reset);
flip_flop16  mod1078(f6PP9,g7PP9,clk,reset);
flip_flop16  mod1079(f6PP10,g7PP10,clk,reset);
flip_flop16  mod1080(f6PP11,g7PP11,clk,reset);
flip_flop16  mod1081(f6PP12,g7PP12,clk,reset);
flip_flop16  mod1082(f6PP13,g7PP13,clk,reset);
flip_flop16  mod1083(f6PP14,g7PP14,clk,reset);
flip_flop16  mod1084(f6PP15,g7PP15,clk,reset);
//FOR STAGE - 8
halfadder mod105(qsum85,qcarry91,carry106,p8);
fulladder mod106(qsum86,qcarry92,g7PP9[0],carry107,sum99);  
fulladder mod107(qsum87,qcarry93,g7PP9[1],carry108,sum100);
fulladder mod108(qsum88,qcarry94,g7PP9[2],carry109,sum101);
fulladder mod109(qsum89,qcarry95,g7PP9[3],carry110,sum102);
fulladder mod110(qsum90,qcarry96,g7PP9[4],carry111,sum103);
fulladder mod111(qsum91,qcarry97,g7PP9[5],carry112,sum104);
fulladder mod112(qsum92,qcarry98,g7PP9[6],carry113,sum105);
fulladder mod113(qsum93,qcarry99,g7PP8[8],carry114,sum106);
fulladder mod114(qsum94,qcarry100,g7PP8[9],carry115,sum107);
fulladder mod115(qsum95,qcarry101,g7PP8[10],carry116,sum108);
fulladder mod116(qsum96,qcarry102,g7PP8[11],carry117,sum109);
fulladder mod117(qsum97,qcarry103,g7PP8[12],carry118,sum110);
fulladder mod118(qsum98,qcarry104,g7PP8[13],carry119,sum111);
fulladder mod119(g7PP7,g7PP8[14],qcarry105,carry120,sum112);
//FOR STAGE - 8 PIPELINE 
flip_flop1  mod479(p07,p08,clk,reset); 
flip_flop1  mod480(p17,p18,clk,reset);
flip_flop1  mod481(p26,p27,clk,reset);
flip_flop1  mod482(p35,p36,clk,reset);
flip_flop1  mod483(p44,p45,clk,reset);
flip_flop1  mod484(p53,p54,clk,reset);
flip_flop1  mod485(p62,p63,clk,reset);
flip_flop1  mod486(p71,p72,clk,reset);
flip_flop1  mod487(p8,p81,clk,reset);
flip_flop1  mod488(carry106,qcarry106,clk,reset); 
flip_flop1  mod489(carry107,qcarry107,clk,reset);
flip_flop1  mod490(carry108,qcarry108,clk,reset);
flip_flop1  mod491(carry109,qcarry109,clk,reset);
flip_flop1  mod492(carry110,qcarry110,clk,reset);
flip_flop1  mod493(carry111,qcarry111,clk,reset);
flip_flop1  mod494(carry112,qcarry112,clk,reset); 
flip_flop1  mod495(carry113,qcarry113,clk,reset); 
flip_flop1  mod496(carry114,qcarry114,clk,reset); 
flip_flop1  mod497(carry115,qcarry115,clk,reset);
flip_flop1  mod498(carry116,qcarry116,clk,reset);
flip_flop1  mod499(carry117,qcarry117,clk,reset);
flip_flop1  mod500(carry118,qcarry118,clk,reset);     
flip_flop1  mod501(carry119,qcarry119,clk,reset);
flip_flop1  mod502(carry120,qcarry120,clk,reset); 
         
flip_flop1  mod503(sum99,qsum99,clk,reset);
flip_flop1  mod504(sum100,qsum100,clk,reset);
flip_flop1  mod505(sum101,qsum101,clk,reset);
flip_flop1  mod506(sum102,qsum102,clk,reset);
flip_flop1  mod507(sum103,qsum103,clk,reset);
flip_flop1  mod508(sum104,qsum104,clk,reset);
flip_flop1  mod509(sum105,qsum105,clk,reset);
flip_flop1  mod510(sum106,qsum106,clk,reset);
flip_flop1  mod511(sum107,qsum107,clk,reset);
flip_flop1  mod512(sum108,qsum108,clk,reset);
flip_flop1  mod513(sum109,qsum109,clk,reset);
flip_flop1  mod514(sum110,qsum110,clk,reset);
flip_flop1  mod515(sum111,qsum111,clk,reset);
flip_flop1  mod516(sum112,qsum112,clk,reset);         
         
flip_flop1 mod1085(g7PP8[15],h8PP8,clk,reset);
flip_flop16  mod1086(g7PP9,h8PP9,clk,reset);
flip_flop16  mod1087(g7PP10,h8PP10,clk,reset);
flip_flop16  mod1088(g7PP11,h8PP11,clk,reset);
flip_flop16  mod1089(g7PP12,h8PP12,clk,reset);
flip_flop16  mod1090(g7PP13,h8PP13,clk,reset);
flip_flop16  mod1091(g7PP14,h8PP14,clk,reset);
flip_flop16  mod1092(g7PP15,h8PP15,clk,reset);
//FOR STAGE - 9
halfadder mod120(qsum99,qcarry106,carry121,p9);
fulladder mod121(qsum100,qcarry107,h8PP10[0],carry122,sum113);  
fulladder mod122(qsum101,qcarry108,h8PP10[1],carry123,sum114);
fulladder mod123(qsum102,qcarry109,h8PP10[2],carry124,sum115);
fulladder mod124(qsum103,qcarry110,h8PP10[3],carry125,sum116);
fulladder mod125(qsum104,qcarry111,h8PP10[4],carry126,sum117);
fulladder mod126(qsum105,qcarry112,h8PP10[5],carry127,sum118);
fulladder mod127(qsum106,qcarry113,h8PP9[7],carry128,sum119);
fulladder mod128(qsum107,qcarry114,h8PP9[8],carry129,sum120);
fulladder mod129(qsum108,qcarry115,h8PP9[9],carry130,sum121);
fulladder mod130(qsum109,qcarry116,h8PP9[10],carry131,sum122);
fulladder mod131(qsum110,qcarry117,h8PP9[11],carry132,sum123);
fulladder mod132(qsum111,qcarry118,h8PP9[12],carry133,sum124);
fulladder mod133(qsum112,qcarry119,h8PP9[13],carry134,sum125);
fulladder mod134(h8PP8,h8PP9[14],qcarry120,carry135,sum126);
//FOR STAGE - 9 PIPELINE 
flip_flop1  mod517(p08,p09,clk,reset); 
flip_flop1  mod518(p18,p19,clk,reset);
flip_flop1  mod519(p27,p28,clk,reset);
flip_flop1  mod520(p36,p37,clk,reset);
flip_flop1  mod521(p45,p46,clk,reset);
flip_flop1  mod522(p54,p55,clk,reset);
flip_flop1  mod523(p63,p64,clk,reset);
flip_flop1  mod524(p72,p73,clk,reset);
flip_flop1  mod525(p81,p82,clk,reset);
flip_flop1  mod526(p9,p91,clk,reset);
flip_flop1  mod527(carry121,qcarry121,clk,reset); 
flip_flop1  mod528(carry122,qcarry122,clk,reset);
flip_flop1  mod529(carry123,qcarry123,clk,reset);
flip_flop1  mod530(carry124,qcarry124,clk,reset);
flip_flop1  mod531(carry125,qcarry125,clk,reset);
flip_flop1  mod532(carry126,qcarry126,clk,reset);
flip_flop1  mod533(carry127,qcarry127,clk,reset); 
flip_flop1  mod534(carry128,qcarry128,clk,reset); 
flip_flop1  mod535(carry129,qcarry129,clk,reset); 
flip_flop1  mod536(carry130,qcarry130,clk,reset);
flip_flop1  mod537(carry131,qcarry131,clk,reset);
flip_flop1  mod538(carry132,qcarry132,clk,reset);
flip_flop1  mod539(carry133,qcarry133,clk,reset);     
flip_flop1  mod540(carry134,qcarry134,clk,reset);
flip_flop1  mod541(carry135,qcarry135,clk,reset); 
         
flip_flop1  mod542(sum113,qsum113,clk,reset);
flip_flop1  mod543(sum114,qsum114,clk,reset);
flip_flop1  mod545(sum115,qsum115,clk,reset);
flip_flop1  mod546(sum116,qsum116,clk,reset);
flip_flop1  mod547(sum117,qsum117,clk,reset);
flip_flop1  mod548(sum118,qsum118,clk,reset);
flip_flop1  mod549(sum119,qsum119,clk,reset);
flip_flop1  mod550(sum120,qsum120,clk,reset);
flip_flop1  mod551(sum121,qsum121,clk,reset);
flip_flop1  mod552(sum122,qsum122,clk,reset);
flip_flop1  mod553(sum123,qsum123,clk,reset);
flip_flop1  mod554(sum124,qsum124,clk,reset);
flip_flop1  mod555(sum125,qsum125,clk,reset);
flip_flop1  mod556(sum126,qsum126,clk,reset);   
   
flip_flop1 mod1093(h8PP9[15],i9PP9,clk,reset);
flip_flop16  mod1094(h8PP10,i9PP10,clk,reset);
flip_flop16  mod1095(h8PP11,i9PP11,clk,reset);
flip_flop16  mod1096(h8PP12,i9PP12,clk,reset);
flip_flop16  mod1097(h8PP13,i9PP13,clk,reset);
flip_flop16  mod1098(h8PP14,i9PP14,clk,reset);
flip_flop16  mod1099(h8PP15,i9PP15,clk,reset); 
//FOR STAGE - 10            
halfadder mod135(qsum113,qcarry121,carry136,p100);
fulladder mod136(qsum114,qcarry122,i9PP11[0],carry137,sum127);  
fulladder mod137(qsum115,qcarry123,i9PP11[1],carry138,sum128);
fulladder mod138(qsum116,qcarry124,i9PP11[2],carry139,sum129);
fulladder mod139(qsum117,qcarry125,i9PP11[3],carry140,sum130);
fulladder mod140(qsum118,qcarry126,i9PP11[4],carry141,sum131);
fulladder mod141(qsum119,qcarry127,i9PP10[6],carry142,sum132);
fulladder mod142(qsum120,qcarry128,i9PP10[7],carry143,sum133);
fulladder mod143(qsum121,qcarry129,i9PP10[8],carry144,sum134);
fulladder mod144(qsum122,qcarry130,i9PP10[9],carry145,sum135);
fulladder mod145(qsum123,qcarry131,i9PP10[10],carry146,sum136);
fulladder mod146(qsum124,qcarry132,i9PP10[11],carry147,sum137);
fulladder mod147(qsum125,qcarry133,i9PP10[12],carry148,sum138);
fulladder mod148(qsum126,qcarry134,i9PP10[13],carry149,sum139);
fulladder mod149(i9PP9,i9PP10[14],qcarry135,carry150,sum140);
//FOR STAGE - 10 PIPELINE 
flip_flop1  mod557(p09,p010,clk,reset); 
flip_flop1  mod558(p19,p110,clk,reset);
flip_flop1  mod559(p28,p29,clk,reset);
flip_flop1  mod560(p37,p38,clk,reset);
flip_flop1  mod561(p46,p47,clk,reset);
flip_flop1  mod562(p55,p56,clk,reset);
flip_flop1  mod563(p64,p65,clk,reset);
flip_flop1  mod564(p73,p74,clk,reset);
flip_flop1  mod565(p82,p83,clk,reset);
flip_flop1  mod566(p91,p92,clk,reset);
flip_flop1  mod567(p100,p101,clk,reset);
flip_flop1  mod568(carry136,qcarry136,clk,reset); 
flip_flop1  mod569(carry137,qcarry137,clk,reset);
flip_flop1  mod570(carry138,qcarry138,clk,reset);
flip_flop1  mod571(carry139,qcarry139,clk,reset);
flip_flop1  mod572(carry140,qcarry140,clk,reset);
flip_flop1  mod573(carry141,qcarry141,clk,reset);
flip_flop1  mod574(carry142,qcarry142,clk,reset); 
flip_flop1  mod575(carry143,qcarry143,clk,reset); 
flip_flop1  mod576(carry144,qcarry144,clk,reset); 
flip_flop1  mod577(carry145,qcarry145,clk,reset);
flip_flop1  mod578(carry146,qcarry146,clk,reset);
flip_flop1  mod579(carry147,qcarry147,clk,reset);
flip_flop1  mod580(carry148,qcarry148,clk,reset);     
flip_flop1  mod581(carry149,qcarry149,clk,reset);
flip_flop1  mod582(carry150,qcarry150,clk,reset); 
         
flip_flop1  mod583(sum127,qsum127,clk,reset);
flip_flop1  mod584(sum128,qsum128,clk,reset);
flip_flop1  mod585(sum129,qsum129,clk,reset);
flip_flop1  mod586(sum130,qsum130,clk,reset);
flip_flop1  mod587(sum131,qsum131,clk,reset);
flip_flop1  mod588(sum132,qsum132,clk,reset);
flip_flop1  mod589(sum133,qsum133,clk,reset);
flip_flop1  mod590(sum134,qsum134,clk,reset);
flip_flop1  mod591(sum135,qsum135,clk,reset);
flip_flop1  mod592(sum136,qsum136,clk,reset);
flip_flop1  mod593(sum137,qsum137,clk,reset);
flip_flop1  mod594(sum138,qsum138,clk,reset);
flip_flop1  mod595(sum139,qsum139,clk,reset);
flip_flop1  mod596(sum140,qsum140,clk,reset);

flip_flop1 mod1200(i9PP10[15],j10PP10,clk,reset);
flip_flop16 mod1100(i9PP11,j10PP11,clk,reset);
flip_flop16 mod1101(i9PP12,j10PP12,clk,reset);
flip_flop16 mod1102(i9PP13,j10PP13,clk,reset);
flip_flop16 mod1103(i9PP14,j10PP14,clk,reset);
flip_flop16 mod1104(i9PP15,j10PP15,clk,reset);
//FOR STAGE - 11
halfadder mod150(qsum127,qcarry136,carry151,p1100);
fulladder mod151(qsum128,qcarry137,j10PP12[0],carry152,sum141);  
fulladder mod152(qsum129,qcarry138,j10PP12[1],carry153,sum142);
fulladder mod153(qsum130,qcarry139,j10PP12[2],carry154,sum143);
fulladder mod154(qsum131,qcarry140,j10PP12[3],carry155,sum144);
fulladder mod155(qsum132,qcarry141,j10PP11[5],carry156,sum145);
fulladder mod156(qsum133,qcarry142,j10PP11[6],carry157,sum146);
fulladder mod240(qsum134,qcarry143,j10PP11[7],carry158,sum147);
fulladder mod157(qsum135,qcarry144,j10PP11[8],carry159,sum148);
fulladder mod158(qsum136,qcarry145,j10PP11[9],carry160,sum149);
fulladder mod159(qsum137,qcarry146,j10PP11[10],carry161,sum150);
fulladder mod160(qsum138,qcarry147,j10PP11[11],carry162,sum151);
fulladder mod161(qsum139,qcarry148,j10PP11[12],carry163,sum152);
fulladder mod162(qsum140,qcarry149,j10PP11[13],carry164,sum153);
fulladder mod163(j10PP10,j10PP11[14],qcarry150,carry165,sum154);
//FOR STAGE - 11 PIPELINE 
flip_flop1  mod597(p010,p011,clk,reset); 
flip_flop1  mod598(p110,p111,clk,reset);
flip_flop1  mod599(p29,p210,clk,reset);
flip_flop1  mod600(p38,p39,clk,reset);
flip_flop1  mod601(p47,p48,clk,reset);
flip_flop1  mod602(p56,p57,clk,reset);
flip_flop1  mod603(p65,p66,clk,reset);
flip_flop1  mod604(p74,p75,clk,reset);
flip_flop1  mod605(p83,p84,clk,reset);
flip_flop1  mod606(p92,p93,clk,reset);
flip_flop1  mod607(p101,p102,clk,reset);
flip_flop1  mod608(p1100,p1101,clk,reset);
flip_flop1  mod609(carry151,qcarry151,clk,reset); 
flip_flop1  mod610(carry152,qcarry152,clk,reset);
flip_flop1  mod611(carry153,qcarry153,clk,reset);
flip_flop1  mod612(carry154,qcarry154,clk,reset);
flip_flop1  mod613(carry155,qcarry155,clk,reset);
flip_flop1  mod614(carry156,qcarry156,clk,reset);
flip_flop1  mod615(carry157,qcarry157,clk,reset); 
flip_flop1  mod616(carry158,qcarry158,clk,reset); 
flip_flop1  mod617(carry159,qcarry159,clk,reset); 
flip_flop1  mod618(carry160,qcarry160,clk,reset);
flip_flop1  mod619(carry161,qcarry161,clk,reset);
flip_flop1  mod620(carry162,qcarry162,clk,reset);
flip_flop1  mod621(carry163,qcarry163,clk,reset);     
flip_flop1  mod622(carry164,qcarry164,clk,reset);
flip_flop1  mod623(carry165,qcarry165,clk,reset); 
         
flip_flop1  mod624(sum141,qsum141,clk,reset);
flip_flop1  mod625(sum142,qsum142,clk,reset);
flip_flop1  mod626(sum143,qsum143,clk,reset);
flip_flop1  mod627(sum144,qsum144,clk,reset);
flip_flop1  mod628(sum145,qsum145,clk,reset);
flip_flop1  mod629(sum146,qsum146,clk,reset);
flip_flop1  mod630(sum147,qsum147,clk,reset);
flip_flop1  mod631(sum148,qsum148,clk,reset);
flip_flop1  mod632(sum149,qsum149,clk,reset);
flip_flop1  mod633(sum150,qsum150,clk,reset);
flip_flop1  mod634(sum151,qsum151,clk,reset);
flip_flop1  mod635(sum152,qsum152,clk,reset);
flip_flop1  mod636(sum153,qsum153,clk,reset);
flip_flop1  mod637(sum154,qsum154,clk,reset);         
         
flip_flop1 mod1105(j10PP11[15],k11PP11,clk,reset);
flip_flop16  mod1106(j10PP12,k11PP12,clk,reset);
flip_flop16  mod1107(j10PP13,k11PP13,clk,reset);
flip_flop16  mod1108(j10PP14,k11PP14,clk,reset);
flip_flop16  mod1109(j10PP15,k11PP15,clk,reset);
//FOR STAGE - 12
halfadder mod164(qsum141,qcarry151,carry166,p1200);
fulladder mod165(qsum142,qcarry152,k11PP13[0],carry167,sum155);  
fulladder mod166(qsum143,qcarry153,k11PP13[1],carry168,sum156);
fulladder mod167(qsum144,qcarry154,k11PP13[2],carry169,sum157);
fulladder mod168(qsum145,qcarry155,k11PP12[4],carry170,sum158);
fulladder mod169(qsum146,qcarry156,k11PP12[5],carry171,sum159);
fulladder mod170(qsum147,qcarry157,k11PP12[6],carry172,sum160);
fulladder mod171(qsum148,qcarry158,k11PP12[7],carry173,sum161);
fulladder mod172(qsum149,qcarry159,k11PP12[8],carry174,sum162);
fulladder mod173(qsum150,qcarry160,k11PP12[9],carry175,sum163);
fulladder mod174(qsum151,qcarry161,k11PP12[10],carry176,sum164);
fulladder mod175(qsum152,qcarry162,k11PP12[11],carry177,sum165);
fulladder mod176(qsum153,qcarry163,k11PP12[12],carry178,sum166);
fulladder mod177(qsum154,qcarry164,k11PP12[13],carry179,sum167);
fulladder mod178(k11PP11,k11PP12[14],qcarry165,carry180,sum168);
//FOR STAGE - 12 PIPELINE 
flip_flop1  mod638(p011,p012,clk,reset); 
flip_flop1  mod639(p111,p112,clk,reset);
flip_flop1  mod640(p210,p211,clk,reset);
flip_flop1  mod641(p39,p310,clk,reset);
flip_flop1  mod642(p48,p49,clk,reset);
flip_flop1  mod643(p57,p58,clk,reset);
flip_flop1  mod644(p66,p67,clk,reset);
flip_flop1  mod645(p75,p76,clk,reset);
flip_flop1  mod646(p84,p85,clk,reset);
flip_flop1  mod647(p93,p94,clk,reset);
flip_flop1  mod648(p102,p103,clk,reset);
flip_flop1  mod649(p1101,p1102,clk,reset);
flip_flop1  mod650(p1200,p1201,clk,reset);
flip_flop1  mod651(carry166,qcarry166,clk,reset); 
flip_flop1  mod652(carry167,qcarry167,clk,reset);
flip_flop1  mod653(carry168,qcarry168,clk,reset);
flip_flop1  mod654(carry169,qcarry169,clk,reset);
flip_flop1  mod655(carry170,qcarry170,clk,reset);
flip_flop1  mod656(carry171,qcarry171,clk,reset);
flip_flop1  mod657(carry172,qcarry172,clk,reset); 
flip_flop1  mod658(carry173,qcarry173,clk,reset); 
flip_flop1  mod659(carry174,qcarry174,clk,reset); 
flip_flop1  mod660(carry175,qcarry175,clk,reset);
flip_flop1  mod661(carry176,qcarry176,clk,reset);
flip_flop1  mod662(carry177,qcarry177,clk,reset);
flip_flop1  mod663(carry178,qcarry178,clk,reset);     
flip_flop1  mod664(carry179,qcarry179,clk,reset);
flip_flop1  mod665(carry180,qcarry180,clk,reset); 
         
flip_flop1  mod666(sum155,qsum155,clk,reset);
flip_flop1  mod667(sum156,qsum156,clk,reset);
flip_flop1  mod668(sum157,qsum157,clk,reset);
flip_flop1  mod669(sum158,qsum158,clk,reset);
flip_flop1  mod670(sum159,qsum159,clk,reset);
flip_flop1  mod671(sum160,qsum160,clk,reset);
flip_flop1  mod672(sum161,qsum161,clk,reset);
flip_flop1  mod673(sum162,qsum162,clk,reset);
flip_flop1  mod674(sum163,qsum163,clk,reset);
flip_flop1  mod675(sum164,qsum164,clk,reset);
flip_flop1  mod676(sum165,qsum165,clk,reset);
flip_flop1  mod677(sum166,qsum166,clk,reset);
flip_flop1  mod678(sum167,qsum167,clk,reset);
flip_flop1  mod679(sum168,qsum168,clk,reset);
         
flip_flop1 mod1110(k11PP12[15],l12PP12,clk,reset);
flip_flop16  mod1111(k11PP13,l12PP13,clk,reset);
flip_flop16  mod1112(k11PP14,l12PP14,clk,reset);
flip_flop16  mod1113(k11PP15,l12PP15,clk,reset);
//FOR STAGE - 13
halfadder mod179(qsum155,qcarry166,carry181,p1300);
fulladder mod180(qsum156,qcarry167,l12PP14[0],carry182,sum169);  
fulladder mod181(qsum157,qcarry168,l12PP14[1],carry183,sum170);
fulladder mod182(qsum158,qcarry169,l12PP13[3],carry184,sum171);
fulladder mod183(qsum159,qcarry170,l12PP13[4],carry185,sum172);
fulladder mod184(qsum160,qcarry171,l12PP13[5],carry186,sum173);
fulladder mod185(qsum161,qcarry172,l12PP13[6],carry187,sum174);
fulladder mod186(qsum162,qcarry173,l12PP13[7],carry188,sum175);
fulladder mod187(qsum163,qcarry174,l12PP13[8],carry189,sum176);
fulladder mod188(qsum164,qcarry175,l12PP13[9],carry190,sum177);
fulladder mod189(qsum165,qcarry176,l12PP13[10],carry191,sum178);
fulladder mod190(qsum166,qcarry177,l12PP13[11],carry192,sum179);
fulladder mod191(qsum167,qcarry178,l12PP13[12],carry193,sum180);
fulladder mod192(qsum168,qcarry179,l12PP13[13],carry194,sum181);
fulladder mod193(l12PP12,l12PP13[14],qcarry180,carry195,sum182);
//FOR STAGE - 13 PIPELINE 
flip_flop1  mod680(p012,p013,clk,reset); 
flip_flop1  mod681(p112,p113,clk,reset);
flip_flop1  mod682(p211,p212,clk,reset);
flip_flop1  mod683(p310,p311,clk,reset);
flip_flop1  mod684(p49,p410,clk,reset);
flip_flop1  mod685(p58,p59,clk,reset);
flip_flop1  mod686(p67,p68,clk,reset);
flip_flop1  mod687(p76,p77,clk,reset);
flip_flop1  mod688(p85,p86,clk,reset);
flip_flop1  mod689(p94,p95,clk,reset);
flip_flop1  mod690(p103,p104,clk,reset);
flip_flop1  mod691(p1102,p1103,clk,reset);
flip_flop1  mod692(p1201,p1202,clk,reset);
flip_flop1  mod693(p1300,p1301,clk,reset);
flip_flop1  mod694(carry181,qcarry181,clk,reset); 
flip_flop1  mod695(carry182,qcarry182,clk,reset);
flip_flop1  mod696(carry183,qcarry183,clk,reset);
flip_flop1  mod697(carry184,qcarry184,clk,reset);
flip_flop1  mod698(carry185,qcarry185,clk,reset);
flip_flop1  mod699(carry186,qcarry186,clk,reset);
flip_flop1  mod700(carry187,qcarry187,clk,reset); 
flip_flop1  mod701(carry188,qcarry188,clk,reset); 
flip_flop1  mod702(carry189,qcarry189,clk,reset); 
flip_flop1  mod703(carry190,qcarry190,clk,reset);
flip_flop1  mod704(carry191,qcarry191,clk,reset);
flip_flop1  mod705(carry192,qcarry192,clk,reset);
flip_flop1  mod706(carry193,qcarry193,clk,reset);     
flip_flop1  mod707(carry194,qcarry194,clk,reset);
flip_flop1  mod708(carry195,qcarry195,clk,reset); 
         
flip_flop1  mod709(sum169,qsum169,clk,reset);
flip_flop1  mod710(sum170,qsum170,clk,reset);
flip_flop1  mod711(sum171,qsum171,clk,reset);
flip_flop1  mod712(sum172,qsum172,clk,reset);
flip_flop1  mod713(sum173,qsum173,clk,reset);
flip_flop1  mod714(sum174,qsum174,clk,reset);
flip_flop1  mod715(sum175,qsum175,clk,reset);
flip_flop1  mod716(sum176,qsum176,clk,reset);
flip_flop1  mod717(sum177,qsum177,clk,reset);
flip_flop1  mod718(sum178,qsum178,clk,reset);
flip_flop1  mod719(sum179,qsum179,clk,reset);
flip_flop1  mod720(sum180,qsum180,clk,reset);
flip_flop1  mod721(sum181,qsum181,clk,reset);
flip_flop1  mod722(sum182,qsum182,clk,reset);   
         
flip_flop1 mod1114(l12PP13[15],m13PP13,clk,reset);
flip_flop16 mod1115(l12PP14,m13PP14,clk,reset);
flip_flop16 mod1116(l12PP15,m13PP15,clk,reset);
//FOR STAGE - 14
halfadder mod194(qsum169,qcarry181,carry196,p1400);
fulladder mod195(qsum170,qcarry182,m13PP15[0],carry197,sum183);  
fulladder mod196(qsum171,qcarry183,m13PP14[2],carry198,sum184);
fulladder mod197(qsum172,qcarry184,m13PP14[3],carry199,sum185);
fulladder mod198(qsum173,qcarry185,m13PP14[4],carry200,sum186);
fulladder mod199(qsum174,qcarry186,m13PP14[5],carry201,sum187);
fulladder mod200(qsum175,qcarry187,m13PP14[6],carry202,sum188);
fulladder mod201(qsum176,qcarry188,m13PP14[7],carry203,sum189);
fulladder mod202(qsum177,qcarry189,m13PP14[8],carry204,sum190);
fulladder mod203(qsum178,qcarry190,m13PP14[9],carry205,sum191);
fulladder mod204(qsum179,qcarry191,m13PP14[10],carry206,sum192);
fulladder mod205(qsum180,qcarry192,m13PP14[11],carry207,sum193);
fulladder mod206(qsum181,qcarry193,m13PP14[12],carry208,sum194);
fulladder mod207(qsum182,qcarry194,m13PP14[13],carry209,sum195);
fulladder mod208(m13PP13,m13PP14[14],qcarry195,carry210,sum196);
//FOR STAGE - 14 PIPELINE 
flip_flop1  mod723(p013,p014,clk,reset); 
flip_flop1  mod724(p113,p114,clk,reset);
flip_flop1  mod725(p212,p213,clk,reset);
flip_flop1  mod726(p311,p312,clk,reset);
flip_flop1  mod727(p410,p411,clk,reset);
flip_flop1  mod728(p59,p510,clk,reset);
flip_flop1  mod729(p68,p69,clk,reset);
flip_flop1  mod730(p77,p78,clk,reset);
flip_flop1  mod731(p86,p87,clk,reset);
flip_flop1  mod732(p95,p96,clk,reset);
flip_flop1  mod733(p104,p105,clk,reset);
flip_flop1  mod734(p1103,p1104,clk,reset);
flip_flop1  mod735(p1202,p1203,clk,reset);
flip_flop1  mod736(p1301,p1302,clk,reset);
flip_flop1  mod737(p1400,p1401,clk,reset);
flip_flop1  mod738(carry196,qcarry196,clk,reset); 
flip_flop1  mod739(carry197,qcarry197,clk,reset);
flip_flop1  mod740(carry198,qcarry198,clk,reset);
flip_flop1  mod741(carry199,qcarry199,clk,reset);
flip_flop1  mod742(carry200,qcarry200,clk,reset);
flip_flop1  mod743(carry201,qcarry201,clk,reset);
flip_flop1  mod744(carry202,qcarry202,clk,reset); 
flip_flop1  mod745(carry203,qcarry203,clk,reset); 
flip_flop1  mod746(carry204,qcarry204,clk,reset); 
flip_flop1  mod747(carry205,qcarry205,clk,reset);
flip_flop1  mod748(carry206,qcarry206,clk,reset);
flip_flop1  mod749(carry207,qcarry207,clk,reset);
flip_flop1  mod750(carry208,qcarry208,clk,reset);     
flip_flop1  mod751(carry209,qcarry209,clk,reset);
flip_flop1  mod752(carry210,qcarry210,clk,reset); 
         
flip_flop1  mod753(sum183,qsum183,clk,reset);
flip_flop1  mod754(sum184,qsum184,clk,reset);
flip_flop1  mod755(sum185,qsum185,clk,reset);
flip_flop1  mod756(sum186,qsum186,clk,reset);
flip_flop1  mod757(sum187,qsum187,clk,reset);
flip_flop1  mod758(sum188,qsum188,clk,reset);
flip_flop1  mod759(sum189,qsum189,clk,reset);
flip_flop1  mod760(sum190,qsum190,clk,reset);
flip_flop1  mod761(sum191,qsum191,clk,reset);
flip_flop1  mod762(sum192,qsum192,clk,reset);
flip_flop1  mod763(sum193,qsum193,clk,reset);
flip_flop1  mod764(sum194,qsum194,clk,reset);
flip_flop1  mod765(sum195,qsum195,clk,reset);
flip_flop1  mod766(sum196,qsum196,clk,reset);
         
flip_flop1 mod1117(m13PP14[15],n14PP14,clk,reset);
flip_flop16 mod1118(m13PP15,n14PP15,clk,reset);
//FOR STAGE - 15
halfadder mod209(qsum183,qcarry196,carry211,p1500);
fulladder mod210(qsum184,qcarry197,n14PP15[1],carry212,sum197);  
fulladder mod211(qsum185,qcarry198,n14PP15[2],carry213,sum198);
fulladder mod212(qsum186,qcarry199,n14PP15[3],carry214,sum199);
fulladder mod213(qsum187,qcarry200,n14PP15[4],carry215,sum200);
fulladder mod214(qsum188,qcarry201,n14PP15[5],carry216,sum201);
fulladder mod215(qsum189,qcarry202,n14PP15[6],carry217,sum202);
fulladder mod216(qsum190,qcarry203,n14PP15[7],carry218,sum203);
fulladder mod217(qsum191,qcarry204,n14PP15[8],carry219,sum204);
fulladder mod218(qsum192,qcarry205,n14PP15[9],carry220,sum205);
fulladder mod219(qsum193,qcarry206,n14PP15[10],carry221,sum206);
fulladder mod220(qsum194,qcarry207,n14PP15[11],carry222,sum207);
fulladder mod221(qsum195,qcarry208,n14PP15[12],carry223,sum208);
fulladder mod222(qsum196,qcarry209,n14PP15[13],carry224,sum209);
fulladder mod223(n14PP14,n14PP15[14],qcarry210,carry225,sum210);
//FOR STAGE - 15 PIPELINE 
flip_flop1  mod767(p014,p015,clk,reset); 
flip_flop1  mod768(p114,p115,clk,reset);
flip_flop1  mod769(p213,p214,clk,reset);
flip_flop1  mod770(p312,p313,clk,reset);
flip_flop1  mod771(p411,p412,clk,reset);
flip_flop1  mod772(p510,p511,clk,reset);
flip_flop1  mod773(p69,p610,clk,reset);
flip_flop1  mod774(p78,p79,clk,reset);
flip_flop1  mod775(p87,p88,clk,reset);
flip_flop1  mod776(p96,p97,clk,reset);
flip_flop1  mod777(p105,p106,clk,reset);
flip_flop1  mod778(p1104,p1105,clk,reset);
flip_flop1  mod779(p1203,p1204,clk,reset);
flip_flop1  mod780(p1302,p1303,clk,reset);
flip_flop1  mod781(p1401,p1402,clk,reset);
flip_flop1  mod782(p1500,p1501,clk,reset);
flip_flop1  mod783(carry211,qcarry211,clk,reset); 
flip_flop1  mod784(carry212,qcarry212,clk,reset);
flip_flop1  mod785(carry213,qcarry213,clk,reset);
flip_flop1  mod786(carry214,qcarry214,clk,reset);
flip_flop1  mod787(carry215,qcarry215,clk,reset);
flip_flop1  mod788(carry216,qcarry216,clk,reset);
flip_flop1  mod789(carry217,qcarry217,clk,reset); 
flip_flop1  mod790(carry218,qcarry218,clk,reset); 
flip_flop1  mod791(carry219,qcarry219,clk,reset); 
flip_flop1  mod792(carry220,qcarry220,clk,reset);
flip_flop1  mod793(carry221,qcarry221,clk,reset);
flip_flop1  mod794(carry222,qcarry222,clk,reset);
flip_flop1  mod795(carry223,qcarry223,clk,reset);     
flip_flop1  mod796(carry224,qcarry224,clk,reset);
flip_flop1  mod797(carry225,qcarry225,clk,reset); 
         
flip_flop1  mod798(sum197,qsum197,clk,reset);
flip_flop1  mod799(sum198,qsum198,clk,reset);
flip_flop1  mod800(sum199,qsum199,clk,reset);
flip_flop1  mod801(sum200,qsum200,clk,reset);
flip_flop1  mod802(sum201,qsum201,clk,reset);
flip_flop1  mod803(sum202,qsum202,clk,reset);
flip_flop1  mod804(sum203,qsum203,clk,reset);
flip_flop1  mod805(sum204,qsum204,clk,reset);
flip_flop1  mod806(sum205,qsum205,clk,reset);
flip_flop1  mod807(sum206,qsum206,clk,reset);
flip_flop1  mod808(sum207,qsum207,clk,reset);
flip_flop1  mod809(sum208,qsum208,clk,reset);
flip_flop1  mod810(sum209,qsum209,clk,reset);
flip_flop1  mod811(sum210,qsum210,clk,reset); 
         
flip_flop1 mod1119(n14PP15[15],o15PP15,clk,reset);
//FOR STAGE - 16
halfadder mod224(qsum197,qcarry211,carry226,p1600);
fulladder mod225(qsum198,qcarry212,carry226,carry227,p1700);  
fulladder mod226(qsum199,qcarry213,carry227,carry228,p1800);
fulladder mod227(qsum200,qcarry214,carry228,carry229,p1900);
fulladder mod228(qsum201,qcarry215,carry229,carry230,p2000);
fulladder mod229(qsum202,qcarry216,carry230,carry231,p2100);
fulladder mod230(qsum203,qcarry217,carry231,carry232,p2200);
fulladder mod231(qsum204,qcarry218,carry232,carry233,p2300);
fulladder mod232(qsum205,qcarry219,carry233,carry234,p2400);
fulladder mod233(qsum206,qcarry220,carry234,carry235,p2500);
fulladder mod234(qsum207,qcarry221,carry235,carry236,p2600);
fulladder mod235(qsum208,qcarry222,carry236,carry237,p2700);
fulladder mod236(qsum209,qcarry223,carry237,carry238,p2800);
fulladder mod237(qsum210,qcarry224,carry238,carry239,p2900);
fulladder mod238(o15PP15,qcarry225,carry239,p3100,p3000);


assign out = {p3100,p3000,p2900,p2800,p2700,p2600,p2500,p2400,p2300,p2200,p2100,p2000,p1900,p1800,p1700,p1600,p1501,p1402,p1303,p1204,p1105,p106,p97,p88,p79,p610,p511,p412,p313,p214,p115,p015};    

endmodule